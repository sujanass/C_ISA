class C_ISA_addi4sp_sequence extends C_ISA_sequence;
//factory registration
`uvm_object_utils(C_ISA_addi4sp_sequence)

  //creating sequence item handle
C_ISA_seq_item seq_item;

int scenario;

//function new constructor
function new(string name="C_ISA_addi4sp_sequence");
super.new(name);
endfunction

//build phase
function build_phase(uvm_phase, phase);
//super.new(phase);
seq_item = C_ISA_seq_item::type_id::create("seq_item");
endfunction

//task
task body();

//reset scenario
`uvm_info (get_type_name(),"addi4sp sequence: inside body", UVM_LOW)

 if (scenario == 1)
       // repeat(5) 
       begin
        `uvm_do_with(seq_item,{
	seq_item.risc_rst        	== 1'b0;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b000;	//rd'+8 
	seq_item.instruction[12:5]      == 8'b00000000;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;		
	});
	
	end

 if (scenario == 2)
   //   repeat(2) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b000;	//rd'+8
	seq_item.instruction[12:5]      == 8'b00000010;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

 if (scenario == 3)
    //  repeat(2) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b010;	//rd'+8
	seq_item.instruction[12:5]      == 8'b00000000;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

  if (scenario == 4)
    //  repeat(2) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b011;	//rd'+8
	seq_item.instruction[12:5]      == 8'b00000011;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

  if (scenario == 5)
  //    repeat(2) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
//	seq_item.instruction[4:2]       == 3'b000;	//rd'+8
	seq_item.instruction[12:5]      == 8'b00000100;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

if (scenario == 6)
    //  repeat(10) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b000;	//rd'+8
	seq_item.instruction[12:5]      == 8'b11111111;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

if (scenario == 7)
     // repeat(2) 
       begin
        `uvm_do_with(seq_item,{
  	seq_item.risc_rst        	== 1'b1;
	seq_item.instruction[1:0]       == 2'b00;	//opcode(00)
	seq_item.instruction[4:2]       == 3'b001;	//rd'+8
	seq_item.instruction[12:5]      == 8'b00000110;	//imm[5:4|9:6|2|3]
	seq_item.instruction[15:13]     == 3'b000;	//funct3(000)
	seq_item.data_mem_read_data_i   == 32'b0;	
	});
	end

endtask

endclass

class C_ISA_all_test extends uvm_test;

  //factory registration
  `uvm_component_utils(C_ISA_all_test)

  //creating environment and sequence handle
  C_ISA_env env;
  C_ISA_all_sequence all_seq;
  
  //constructor
  function new(string name = "C_ISA_all_test",uvm_component parent=null);
    super.new(name,parent);
  endfunction
 
  //build phase
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = C_ISA_env::type_id::create("env",this); 
    all_seq = C_ISA_all_sequence::type_id::create("all_seq"); 
  endfunction


//end of elaboration phase
	function void end_of_elaboration_phase(uvm_phase phase);
		uvm_top.print_topology();
	endfunction

task run_phase(uvm_phase phase);
    phase.raise_objection(this);
  //  #100;
   `uvm_info(get_name(),$sformatf("inside the base all_test"),UVM_MEDIUM)

   begin
all_seq.scenario = 1;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 1 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 2;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 2 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 3;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 3 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 4;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 4 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 5;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 5 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 6;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 6 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 7;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 7 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 8;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 8 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 9;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 9 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 10;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 10 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 11;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 11 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 12;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 12 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 13;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 13 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 14;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 14 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 15;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 15 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 16;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 16 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 17;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 17 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 18;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 18 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 19;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 19 is completed"),UVM_MEDIUM)
end

begin
all_seq.scenario = 20;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 20 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 21;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 21 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 22;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 22 is completed"),UVM_MEDIUM)
end 

begin
all_seq.scenario = 23;
all_seq.start(env.agent.sequencer);
`uvm_info(get_type_name(),$sformatf("all_test scenario 23 is completed"),UVM_MEDIUM)
end 

    phase.drop_objection(this);

	phase.phase_done.set_drain_time(this,100);
   
  endtask

endclass 

